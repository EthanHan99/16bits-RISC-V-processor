library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

-----------Entity Declaration----------------------------
entity DMEM is
  port( Rls : in std_logic_vector(7 downto 0);
    Ry : in std_logic_vector(7 downto 0);
    Reg_Ind : in std_logic;
    ALUop : in std_logic_vector(3 downto 0);
    memd : in std_logic_vector(7 downto 0);
    MEM_op : out std_logic_vector(7 downto 0));
  end entity DMEM;
-----------------------------------------------------------
  
----------------------------Architecture Body Declaration------------------------------------------------------------------------
  architecture DMEM_arch of DMEM is
    signal daddr : std_logic_vector(7 downto 0);
  
    -------Componet Declaration--------------------    
    component MUX2_1 is
     port( Ry : in std_logic_vector(7 downto 0);
      IM : in std_logic_vector(7 downto 0);
      SEL : in std_logic;
      To_ALU : out std_logic_vector(7 downto 0));
    end component MUX2_1;
    ----------------------------------------------- 
      
            
    begin     --architecture begins here
      --------Port Map----------------------
      MUX1 : MUX2_1 port map(
                      Ry => Rls,
                      IM => Ry,
                      SEL => Reg_Ind,
                      To_ALU => daddr);
      ----------------------------------------                       
                      
      ---------------Process------------------------------------------------------------------------------------------------------------                
      PMUX1 : process(daddr)
      type DMEM_array is array(255 downto 0) of std_logic_vector(7 downto 0);
      variable data_mem_array : DMEM_array := ("00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","00000000","00000000","00000000","00000000","00000000",
                                            "00000000","00000000","00000000","10101010","11110000","00001111","11001100","00110011");
                                                                 
      
      begin     --Process begins here
        case ALUop(3 downto 0)  is
        when "1000" => MEM_op <=  data_mem_array(conv_integer(daddr));
        when "1001" => data_mem_array(conv_integer(memd)) := daddr;
        when "1010" => MEM_op <= data_mem_array(conv_integer(daddr));
        when "1011" => data_mem_array(conv_integer(daddr)) := memd;
        when  others => null;
      end case;
    end process PMUX1; --Process ends here
                            
end architecture DMEM_arch;     --architecture ends here 